module demultiplexer(d,s,y);
input d;
input [2:0]s;
output [7:0]y;
endmodule
